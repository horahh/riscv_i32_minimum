module alu_connections(
   wire clock,
   wirte enable,
